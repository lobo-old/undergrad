library verilog;
use verilog.vl_types.all;
entity bascule_vlg_vec_tst is
end bascule_vlg_vec_tst;
