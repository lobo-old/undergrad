library verilog;
use verilog.vl_types.all;
entity BLOCK2_vlg_vec_tst is
end BLOCK2_vlg_vec_tst;
