library verilog;
use verilog.vl_types.all;
entity tuto_vlg_sample_tst is
    port(
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end tuto_vlg_sample_tst;
