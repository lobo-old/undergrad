library verilog;
use verilog.vl_types.all;
entity test_Tog_flipflop_vlg_vec_tst is
end test_Tog_flipflop_vlg_vec_tst;
