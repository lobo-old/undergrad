library verilog;
use verilog.vl_types.all;
entity tuto_vlg_vec_tst is
end tuto_vlg_vec_tst;
