library verilog;
use verilog.vl_types.all;
entity compteurModule10_vlg_vec_tst is
end compteurModule10_vlg_vec_tst;
