library verilog;
use verilog.vl_types.all;
entity SCOMP2_vlg_vec_tst is
end SCOMP2_vlg_vec_tst;
