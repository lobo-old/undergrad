library verilog;
use verilog.vl_types.all;
entity adicionaire1_vlg_vec_tst is
end adicionaire1_vlg_vec_tst;
