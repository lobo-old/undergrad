library verilog;
use verilog.vl_types.all;
entity CompteurN_vlg_vec_tst is
end CompteurN_vlg_vec_tst;
