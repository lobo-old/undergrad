library verilog;
use verilog.vl_types.all;
entity Compteur16_vlg_vec_tst is
end Compteur16_vlg_vec_tst;
