library verilog;
use verilog.vl_types.all;
entity adicionaire1 is
    port(
        r               : out    vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        s               : out    vl_logic
    );
end adicionaire1;
