library verilog;
use verilog.vl_types.all;
entity test_TFF_vlg_vec_tst is
end test_TFF_vlg_vec_tst;
