library verilog;
use verilog.vl_types.all;
entity compteur4bits_vlg_vec_tst is
end compteur4bits_vlg_vec_tst;
