library verilog;
use verilog.vl_types.all;
entity adicionaire1BIT_vlg_vec_tst is
end adicionaire1BIT_vlg_vec_tst;
