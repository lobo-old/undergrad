library verilog;
use verilog.vl_types.all;
entity adicionaire1BIT_vlg_check_tst is
    port(
        r               : in     vl_logic;
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end adicionaire1BIT_vlg_check_tst;
